/*

Copyright (c) 2016 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * Testbench for lfsr
 */
module test_lfsr_prbs9;

// Parameters
parameter LFSR_WIDTH = 9;
parameter LFSR_POLY = 9'h021;
parameter LFSR_CONFIG = "FIBONACCI";
parameter LFSR_FEED_FORWARD = 0;
parameter REVERSE = 0;
parameter DATA_WIDTH = 8;
parameter STYLE = "AUTO";

// Inputs
reg clk = 0;
reg rst = 0;
reg [7:0] current_test = 0;

reg [DATA_WIDTH-1:0] data_in = 0;
reg [LFSR_WIDTH-1:0] state_in = 0;

// Outputs
wire [DATA_WIDTH-1:0] data_out;
wire [LFSR_WIDTH-1:0] state_out;

initial begin
    // myhdl integration
    $from_myhdl(
        clk,
        rst,
        current_test,
        data_in,
        state_in
    );
    $to_myhdl(
        data_out,
        state_out
    );

    // dump file
    $dumpfile("test_lfsr_prbs9.lxt");
    $dumpvars(0, test_lfsr_prbs9);
end

lfsr #(
    .LFSR_WIDTH(LFSR_WIDTH),
    .LFSR_POLY(LFSR_POLY),
    .LFSR_CONFIG(LFSR_CONFIG),
    .LFSR_FEED_FORWARD(LFSR_FEED_FORWARD),
    .REVERSE(REVERSE),
    .DATA_WIDTH(DATA_WIDTH),
    .STYLE(STYLE)
)
UUT (
    .data_in(data_in),
    .state_in(state_in),
    .data_out(data_out),
    .state_out(state_out)
);

endmodule
